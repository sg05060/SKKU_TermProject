module Controller(
    
)