module Custom_Addr_Decoder(
    input [4:0] cnt,            // stage 27 -> 2^5 = 32
    output reg [5:0] addr       // 
);
    always @(*) begin
        case(cnt)
            5'b0_0000 : addr = 6'b00_0000;
            5'b0_0001 : addr = 6'b00_0001;
            5'b0_0010 : addr = 6'b00_0010;
            5'b0_0011 : addr = 6'b00_0011;
            5'b0_0100 : addr = 6'b00_1001;
            5'b0_0101 : addr = 6'b00_1010;
            5'b0_0110 : addr = 6'b00_1011;
            5'b0_0111 : addr = 6'b00_1100;
            5'b0_1000 : addr = 6'b00_1101;
            5'b0_1001 : addr = 6'b00_1110;
            5'b0_1010 : addr = 6'b00_0100;
            5'b0_1011 : addr = 6'b00_1111;
            5'b0_1100 : addr = 6'b00_0101;
            5'b0_1101 : addr = 6'b01_0000;
            5'b0_1110 : addr = 6'b00_0110;
            5'b0_1111 : addr = 6'b01_0001;
            5'b1_0000 : addr = 6'b01_0010;
            5'b1_0001 : addr = 6'b00_0111;
            5'b1_0010 : addr = 6'b01_0011;
            5'b1_0011 : addr = 6'b00_1000;
            5'b1_0100 : addr = 6'b01_0100;
            5'b1_0101 : addr = 6'b01_0101;
            5'b1_0110 : addr = 6'b01_0110;
            5'b1_0111 : addr = 6'b01_0111;
            5'b1_1000 : addr = 6'b01_1000;
            default   : addr = 6'b00_0000;
        endcase
    end
    
    // binary output expression
    // 11000 011000
    // 10010 000001
    // 10011 001000
    // 10001 000110
    // 01-00 000001
    // 011-1 010000
    // 0100- 001000
    // 00111 001100
    // 00101 001010
    // 0-110 000010
    // 01-11 000001
    // 1011- 000010
    // -0001 000001
    // 101-1 000001
    // 100-0 010010
    // 01--0 000100
    // 001-0 001001
    // 0-011 000011
    // -0-10 000010
    // 010-1 001110
    // 101-- 010100
    
    // boolean expression
    // addr[5] = none
    // addr[4] = 11000 | 011-1 | 100-0 | 101--
    // addr[3] = 11000 | 10011 | 0100- | 00111 | 00101 | 001-0 | 010-1
    // addr[2] = 10001 | 00111 | 01--0 | 010-1 | 101--
    // addr[1] = 10001 | 00101 | 0-110 | 1011- | 100-0 | 0-011 | -0-10 | 010-1
    // addr[0] = 10010 | 01-00 | 01-11 | -0001 | 101-1 | 001-0 | 0-011

endmodule