module Custom_ACC_en_Decoder(
    input [4:0] cnt,            // stage 27 -> 2^5 = 32
    output reg [3:0] acc_en     // 
);
    always @(*) begin
        case(cnt)
            5'b0_0000 : acc_en = 4'b0000;
            5'b0_0001 : acc_en = 4'b0000;
            5'b0_0010 : acc_en = 4'b0000;
            5'b0_0011 : acc_en = 4'b0000;
            5'b0_0100 : acc_en = 4'b0000;
            5'b0_0101 : acc_en = 4'b1000;
            5'b0_0110 : acc_en = 4'b1100;
            5'b0_0111 : acc_en = 4'b1100;
            5'b0_1000 : acc_en = 4'b0100;
            5'b0_1001 : acc_en = 4'b1010;
            5'b0_1010 : acc_en = 4'b0111;
            5'b0_1011 : acc_en = 4'b1000;
            5'b0_1100 : acc_en = 4'b0111;
            5'b0_1101 : acc_en = 4'b1000;
            5'b0_1110 : acc_en = 4'b0101;
            5'b0_1111 : acc_en = 4'b0000;
            5'b1_0000 : acc_en = 4'b1010;
            5'b1_0001 : acc_en = 4'b0111;
            5'b1_0010 : acc_en = 4'b1000;
            5'b1_0011 : acc_en = 4'b0111;
            5'b1_0100 : acc_en = 4'b1000;
            5'b1_0101 : acc_en = 4'b0101;
            5'b1_0110 : acc_en = 4'b0010;
            5'b1_0111 : acc_en = 4'b0011;
            5'b1_1000 : acc_en = 4'b0011;
            5'b1_1001 : acc_en = 4'b0001;
            default   : acc_en = 4'b0000;
        endcase
    end
    
    // binary output expression
    // 01010 0010
    // 01001 0010
    // 01100 0011
    // 01-10 0001
    // 0-101 1000
    // 1011- 0010
    // 0011- 1100
    // 11000 0011
    // 010-1 1000
    // 10-01 0100
    // 10-00 1000
    // 100-0 1000
    // 1-001 0001
    // 1000- 0010
    // 01--0 0100
    // 100-1 0110
    // 10--1 0001
    
    // Boolean expression of acc_en[3:0]
    // acc_en[3] = 0-101 | 0011- | 010-1 | 10-00 | 100-0
    // acc_en[2] = 0011- | 10-01 | 01--0 | 100-1
    // acc_en[1] = 01010 | 01001 | 01100 | 1011- | 11000 | 1000- | 100-1
    // acc_en[0] = 01100 | 01-10 | 11000 | 1-001 | 10--1
    
    
endmodule